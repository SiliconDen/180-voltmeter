.ALIAS cap_mim_2f0ff mim_2p0fF
.end
