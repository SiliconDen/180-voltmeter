.ALIAS cap_mim_2f0fF mim_2p0ff
